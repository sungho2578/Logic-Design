`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   09:26:08 11/08/2018
// Design Name:   EdgeDetector
// Module Name:   C:/Users/SH-HP/UCR/CS 120A/Lab4/Lab4_Part2/EdgeDetectorTb.v
// Project Name:  Lab4_Part2
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: EdgeDetector
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module EdgeDetectorTb;

	// Outputs
	wire ;

	// Instantiate the Unit Under Test (UUT)
	EdgeDetector uut (
		.()
	);

	initial begin
		// Initialize Inputs

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

